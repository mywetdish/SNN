interface in_intf(input logic clk, input logic rst);

    bit [961-1:0] spike_i;

endinterface