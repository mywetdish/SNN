class out_transaction;
    logic [2:0] spike_o;
endclass