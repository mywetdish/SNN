class in_transaction;
    bit [961-1:0] spike_i;

    //constraint c_spike { spike_i < 1024*1024; }
endclass