interface out_intf(input logic clk, input logic rst);
    bit [2:0] spike_o;
    bit       valid_spike;
endinterface